package Types;
typedef logic [REG_WIDTH-1:0] register;
typedef logic [INSTR_WIDTH-1:0] instr;
endpackage: Types

